
`timescale   1ns/1ps
//--------------------------------------------------------------------------------------------------
// interface def
//--------------------------------------------------------------------------------------------------
interface apb3_if 
#(
	parameter DW = 32,	
	parameter AW = 32
)(
	input clk,
	input rstn
);	
	//----------------------------------------------------------------------------------------------
	// logic define
	//----------------------------------------------------------------------------------------------
	logic 	[AW - 1 : 0]	addr;  
	logic 					enable;
	logic 	[DW - 1 : 0]	rdata; 
	logic 					ready; 
	logic 					sel;  
	logic 					slverr;
	logic 	[DW - 1 : 0]	wdata; 
	logic 					write;
	
	//----------------------------------------------------------------------------------------------
	// modport define
	//----------------------------------------------------------------------------------------------	
	modport m (
		input 	clk, rstn,
		output	addr, enable, sel, wdata, write,
		input 	rdata, ready, slverr
	);
	
	modport s (
		input 	clk, rstn,
		input	addr, enable, sel, wdata, write,
		output 	rdata, ready, slverr
	);

endinterface
//--------------------------------------------------------------------------------------------------
// eof
//--------------------------------------------------------------------------------------------------

